library verilog;
use verilog.vl_types.all;
entity decoder7_vlg_vec_tst is
end decoder7_vlg_vec_tst;
